module ID_stage (
    input clk,    // Clock
    input rst  // Asynchronous reset active high
    // input [31:0] Instruction,
    // output [31:0] reg1, reg2,
    // input [4:0] src1, src2
    // output IF_flush,
    // output [4:0] Dest,
    // output [31:0] Reg2, Val2, Val1,
    // output Br_taken,
    // output [3:0] EXE_CMD,
    // output MEM_R_EN, MEM_W_EN, WB_EN
);

// Register_file register_file(clk, rst, src1, src2, reg1, reg2);


endmodule