module Control_unit (
    input clk,    // Clock
    input rst  // Asynchronous reset active low
);

endmodule